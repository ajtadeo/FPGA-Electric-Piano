module piano
  (
    clk,
    SW_C, SW_D, SW_E, SW_F, SW_G, SW_A, SW_B,
    BTN_R, BTN_L, BTN_U, BTN_D
  );

  input clk;

  input SW_C;
  input SW_D;
  input SW_E;
  input SW_F;
  input SW_G;
  input SW_A;
  input SW_B;

  input BTN_R;
  input BTN_L;
  input BTN_U;
  input BTN_D;

  wire clk_1;
  wire clk_2;
  wire clk_4;
  wire clk_256;

  clocks clks(.clk_100M(clk),
    .clk_1(clk_1), .clk_2(clk_2), .clk_4(clk_4), .clk_256(clk_256)
  );

  wire rst;
  wire [6:0] note_switches;
  wire toggle_pb;
  wire inc_octave;
  wire dec_octave;

  debounced inputs(.clk(clk_256),
    .SW_C(SW_C),
    .SW_D(SW_D),
    .SW_E(SW_E),
    .SW_F(SW_F),
    .SW_G(SW_G),
    .SW_A(SW_A),
    .SW_B(SW_B),
    .BTN_R(BTN_R), .BTN_R(BTN_L),
    .BTN_R(BTN_U), .BTN_R(BTN_D),
    .note_switches(note_switches),
    .rst(rst), .toggle_pb(toggle_pb),
    .inc_octave(inc_octave), .dec_octave(dec_octave)
  );

  always @ (posedge ^note_switches or posedge ~^note_switches) begin
    if (!pb_mode) begin
      // DO STUFF
    end
  end
endmodule
